-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Jun 18 09:57:11 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Controller IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        go : IN STD_LOGIC := '0';
        NZ : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        code : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
        choice : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        load_AC : OUT STD_LOGIC;
        load_PC : OUT STD_LOGIC;
        load_REM : OUT STD_LOGIC;
        load_RDM : OUT STD_LOGIC;
        load_RI : OUT STD_LOGIC;
        load_NZ : OUT STD_LOGIC;
        selREM : OUT STD_LOGIC;
        selRDM : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        selUAL : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        sumPC : OUT STD_LOGIC;
        writeOn : OUT STD_LOGIC;
        readOn : OUT STD_LOGIC;
        turnDspOn : OUT STD_LOGIC
    );
END Controller;

ARCHITECTURE BEHAVIOR OF Controller IS
    TYPE type_fstate IS (Search2,Search1,Search3,Check,NOP,NOT1,PREP2,PREP3,PREP1,STA1,STA2,PREP4,LDA,AND1,OR1,ADD,HLT,JnNZ,JZ,JMP3,JMP2,JMP1,JN,SetAdress1,SetData,Decision,Wait1,LoadAC,Start,DISP1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,go,NZ,code,choice)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Start;
            load_AC <= '0';
            load_PC <= '0';
            load_REM <= '0';
            load_RDM <= '0';
            load_RI <= '0';
            load_NZ <= '0';
            selREM <= '0';
            selRDM <= "00";
            selUAL <= "000";
            sumPC <= '0';
            writeOn <= '0';
            readOn <= '0';
            turnDspOn <= '0';
        ELSE
            load_AC <= '0';
            load_PC <= '0';
            load_REM <= '0';
            load_RDM <= '0';
            load_RI <= '0';
            load_NZ <= '0';
            selREM <= '0';
            selRDM <= "00";
            selUAL <= "000";
            sumPC <= '0';
            writeOn <= '0';
            readOn <= '0';
            turnDspOn <= '0';
            CASE fstate IS
                WHEN Search2 =>
                    reg_fstate <= Search3;

                    sumPC <= '1';

                    load_RDM <= '1';

                    readOn <= '1';

                    selRDM <= "00";
                WHEN Search1 =>
                    reg_fstate <= Search2;

                    load_REM <= '1';

                    selREM <= '0';
                WHEN Search3 =>
                    IF ((go = '1')) THEN
                        reg_fstate <= Check;
                    ELSIF ((go = '0')) THEN
                        reg_fstate <= Search3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Search3;
                    END IF;

                    load_RI <= '1';

                    readOn <= '1';

                    turnDspOn <= '1';
                WHEN Check =>
                    IF ((code(3 DOWNTO 0) = "0110")) THEN
                        reg_fstate <= NOT1;
                    ELSIF ((((((code(3 DOWNTO 0) = "0001") OR (code(3 DOWNTO 0) = "0010")) OR (code(3 DOWNTO 0) = "0011")) OR (code(3 DOWNTO 0) = "0100")) OR (code(3 DOWNTO 0) = "0101"))) THEN
                        reg_fstate <= PREP1;
                    ELSIF ((code(3 DOWNTO 0) = "1001")) THEN
                        reg_fstate <= JZ;
                    ELSIF ((code(3 DOWNTO 0) = "1010")) THEN
                        reg_fstate <= JN;
                    ELSIF ((code(3 DOWNTO 0) = "1111")) THEN
                        reg_fstate <= HLT;
                    ELSIF ((code(3 DOWNTO 0) = "1000")) THEN
                        reg_fstate <= JMP1;
                    ELSE
                        reg_fstate <= NOP;
                    END IF;
                WHEN NOP =>
                    reg_fstate <= Wait1;
                WHEN NOT1 =>
                    reg_fstate <= Wait1;

                    selUAL <= "011";

                    load_AC <= '1';
                WHEN PREP2 =>
                    reg_fstate <= PREP3;

                    sumPC <= '1';

                    load_RDM <= '1';

                    readOn <= '1';

                    selRDM <= "00";
                WHEN PREP3 =>
                    IF ((code(3 DOWNTO 0) = "0001")) THEN
                        reg_fstate <= STA1;
                    ELSE
                        reg_fstate <= PREP4;
                    END IF;

                    load_REM <= '1';

                    selREM <= '1';
                WHEN PREP1 =>
                    reg_fstate <= PREP2;

                    load_REM <= '1';

                    selREM <= '0';
                WHEN STA1 =>
                    reg_fstate <= STA2;

                    load_RDM <= '1';

                    selRDM <= "01";
                WHEN STA2 =>
                    reg_fstate <= Wait1;

                    writeOn <= '1';
                WHEN PREP4 =>
                    IF ((code(3 DOWNTO 0) = "0010")) THEN
                        reg_fstate <= LDA;
                    ELSIF ((code(3 DOWNTO 0) = "0011")) THEN
                        reg_fstate <= ADD;
                    ELSIF ((code(3 DOWNTO 0) = "0100")) THEN
                        reg_fstate <= AND1;
                    ELSIF ((code(3 DOWNTO 0) = "0101")) THEN
                        reg_fstate <= OR1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= PREP4;
                    END IF;

                    load_RDM <= '1';

                    readOn <= '1';

                    selRDM <= "00";
                WHEN LDA =>
                    reg_fstate <= Wait1;

                    selUAL <= "100";

                    load_AC <= '1';

                    load_NZ <= '1';
                WHEN AND1 =>
                    reg_fstate <= Wait1;

                    selUAL <= "001";

                    load_AC <= '1';

                    load_NZ <= '1';
                WHEN OR1 =>
                    reg_fstate <= Wait1;

                    selUAL <= "010";

                    load_AC <= '1';

                    load_NZ <= '1';
                WHEN ADD =>
                    reg_fstate <= Wait1;

                    selUAL <= "000";

                    load_AC <= '1';

                    load_NZ <= '1';
                WHEN HLT =>
                    reg_fstate <= HLT;

                    load_REM <= '1';

                    load_RDM <= '1';

                    readOn <= '1';

                    selREM <= '1';

                    selRDM <= "10";

                    turnDspOn <= '1';
                WHEN JnNZ =>
                    reg_fstate <= Wait1;

                    sumPC <= '1';
                WHEN JZ =>
                    IF ((NZ(0) = '0')) THEN
                        reg_fstate <= JnNZ;
                    ELSIF ((NZ(0) = '1')) THEN
                        reg_fstate <= JMP1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= JZ;
                    END IF;
                WHEN JMP3 =>
                    reg_fstate <= Wait1;

                    load_PC <= '1';
                WHEN JMP2 =>
                    reg_fstate <= JMP3;

                    load_RDM <= '1';

                    readOn <= '1';

                    selRDM <= "00";
                WHEN JMP1 =>
                    reg_fstate <= JMP2;

                    load_REM <= '1';

                    selREM <= '0';
                WHEN JN =>
                    IF ((NZ(1) = '1')) THEN
                        reg_fstate <= JMP1;
                    ELSIF ((NZ(1) = '0')) THEN
                        reg_fstate <= JnNZ;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= JN;
                    END IF;
                WHEN SetAdress1 =>
                    IF ((go = '1')) THEN
                        reg_fstate <= SetData;
                    ELSIF ((go = '0')) THEN
                        reg_fstate <= SetAdress1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SetAdress1;
                    END IF;

                    load_REM <= '1';

                    load_RDM <= '1';

                    readOn <= '0';

                    selREM <= '1';

                    selRDM <= "10";

                    turnDspOn <= '1';
                WHEN SetData =>
                    IF ((go = '0')) THEN
                        reg_fstate <= DISP1;
                    ELSIF ((go = '1')) THEN
                        reg_fstate <= SetData;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SetData;
                    END IF;

                    load_RDM <= '1';

                    readOn <= '1';

                    selRDM <= "10";

                    turnDspOn <= '1';

                    writeOn <= '1';
                WHEN Decision =>
                    IF ((choice(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= SetAdress1;
                    ELSIF ((choice(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= Wait1;
                    ELSIF ((choice(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= Decision;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Decision;
                    END IF;
                WHEN Wait1 =>
                    IF ((go = '0')) THEN
                        reg_fstate <= Search1;
                    ELSIF ((go = '1')) THEN
                        reg_fstate <= Wait1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Wait1;
                    END IF;

                    readOn <= '1';

                    turnDspOn <= '1';
                WHEN LoadAC =>
                    IF ((go = '0')) THEN
                        reg_fstate <= Decision;
                    ELSIF ((go = '1')) THEN
                        reg_fstate <= LoadAC;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= LoadAC;
                    END IF;

                    selUAL <= "100";

                    load_AC <= '1';

                    load_RDM <= '1';

                    selRDM <= "10";

                    turnDspOn <= '1';
                WHEN Start =>
                    IF ((go = '1')) THEN
                        reg_fstate <= LoadAC;
                    ELSIF ((go = '0')) THEN
                        reg_fstate <= Start;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Start;
                    END IF;

                    turnDspOn <= '1';
                WHEN DISP1 =>
                    IF ((go = '1')) THEN
                        reg_fstate <= Decision;
                    ELSIF ((go = '0')) THEN
                        reg_fstate <= DISP1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DISP1;
                    END IF;

                    readOn <= '1';

                    turnDspOn <= '1';
                WHEN OTHERS => 
                    load_AC <= 'X';
                    load_PC <= 'X';
                    load_REM <= 'X';
                    load_RDM <= 'X';
                    load_RI <= 'X';
                    load_NZ <= 'X';
                    selREM <= 'X';
                    selRDM <= "XX";
                    selUAL <= "XXX";
                    sumPC <= 'X';
                    writeOn <= 'X';
                    readOn <= 'X';
                    turnDspOn <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
