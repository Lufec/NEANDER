library verilog;
use verilog.vl_types.all;
entity memRAM_vlg_vec_tst is
end memRAM_vlg_vec_tst;
